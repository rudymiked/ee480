##################################################################
##
## Michael Rudy & Russell Brooks
## University of Kentucky
## EE 480 Spring 2014
##
## Module: ROM_ROM_straight.v 
## Dependencies: N/A
##
## Description: initial RAM module for ROM_straight.v program
##
## Last Modified: Michael - 4/24/2014
##
##################################################################
